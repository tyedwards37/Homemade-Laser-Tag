PK   ���WE�t�  Q*     cirkitFile.json�Z�n�F���D{��I[�h�p�>X�$�Q�T)*Nj��;KѺX��d�6d��3ggg�\H�.h�'['Y���mWeS3��`a���쏢0X�u�5���,���]Gݗ����f�Զ��,K3a�E�ͣ4�(�X(�i�	�̮��oV�~��O*#���[D,+X��1�%��"/��({�L�g>�cù���O]��+?u�IV_�{�O�gH;�w�lm������X��41.�x����-bư��0S,b2UQ�i)a�\��%�x|�zϷ�m�Ϛ�i=�}��_�WΟ ��(!!=P�$�0��-B�z��Il���IP�$(z�MD�i؋�40/�wdb� �#s�q=2�>����w�}���3��MƵ]w��<��?
��N��&Aᓠ�IP�$(j=�&"�4������߱���eόM��(/�et2�G��$��~�6}qR柃	�۲��dY���	���-t�W>w>'p��5�0������i>�;L���ܣ\����͍��z��Ӵ�����{�E���e��$�=������˳-�1���=;s�����W��ڗ]����g_� �����Szl��c���]�}�7����+s�Wp��Cv���_]��v��[��ݝ*xk'�:I�D���Ǹ�xP�ǝ�{���l����]�yhxt�^�@�:�c�z=
�*�;u���Lj+�c����y���~
;���J�֚<m��C[T4IU�:�Cl� )��)��T�H�E8-�-2��NA��o�6!��2\�1�T��C�X�z����Mg`��h��m���p��݇s!lfյe�6Z�w�f�������.�u	+�m�hn�կ4��ZY�\��C�*��n�Z���Ghe:�������dݺ��s�����)7E�.���:_;؉�U�L�*��wѫ�"-�b�Õ
���Pp�3�4��,����(����G� �B�d`�����FgT�	�6VCs���0��mV��4�F&c�O錄Ζ�2���C"Y��f1V��+��#b!�©G��>���W�n��	�CX�zXX�Q���� ��1��jI8ߨl͡B�a,�LĔ���WZ�XcE�Y0�""���~�R$�F0�c)�Pz0��3k7�Fa�<ƒs��!��=
��0�/(uK�v�@N9z���L���1�1�H�V2&K��(ч��=l~R��a��1���Yv��:/���8�1�����/�o8��ٛ_/��@��og��Il�gT�j�6�Ґi�vA��JqQZDJ�<"�B&�VFRr[�Z����?"�'���B&��� T:!�;�SN��x�o��hGb�`�:1%�������A��!d�}
��T�,º�"�s��H�Sd!es������*��"�E����u'ͺ��#��T� ��ʾ���8�Y��Ly�p�)c[~\8I�(����X�����M����m{t�ڮ�򡴷�GY�-���#�y0�?��4�9�´�EY����7w�=����F5�=Tkn/�4�~�κeS�݅�=��|>\7���p�}�������=�.	�h��N <%EY�N�"|O
S��B"��WH����R����(wH���S�OG61}��a�D~@�2����g�H)���bx��>�"fP��c���Hm����F��Ԇ�.�U��xk:ۖP� e�W�E����B�3ի�漳7�y�OC��?PK   ���WE�t�  Q*             ��    cirkitFile.jsonPK      =       